module sinWaveGenerator(
	input CLK,
	output signed [15:0] sinOut
	);
	
	logic [31:0] x = 0;
	
	logic CLK_Sin = 0;
	logic [31:0] counter = 0;
	
	logic signed [31:0] sin = 0;
	
	assign sinOut = sin[15:0];
	
	always @(posedge CLK)begin
		if(counter < 111)begin
			counter <= counter + 1;
		end
		else begin
			counter <= 0;
			CLK_Sin <= ~CLK_Sin;
		end
	end
	
	always @(posedge CLK_Sin)begin
		case(x)
			0 : sin <= 0;
			1 : sin <= 6;
			2 : sin <= 13;
			3 : sin <= 19;
			4 : sin <= 25;
			5 : sin <= 31;
			6 : sin <= 38;
			7 : sin <= 44;
			8 : sin <= 50;
			9 : sin <= 56;
			10 : sin <= 62;
			11 : sin <= 68;
			12 : sin <= 74;
			13 : sin <= 80;
			14 : sin <= 86;
			15 : sin <= 92;
			16 : sin <= 98;
			17 : sin <= 104;
			18 : sin <= 109;
			19 : sin <= 115;
			20 : sin <= 121;
			21 : sin <= 126;
			22 : sin <= 132;
			23 : sin <= 137;
			24 : sin <= 142;
			25 : sin <= 147;
			26 : sin <= 152;
			27 : sin <= 157;
			28 : sin <= 162;
			29 : sin <= 167;
			30 : sin <= 172;
			31 : sin <= 177;
			32 : sin <= 181;
			33 : sin <= 185;
			34 : sin <= 190;
			35 : sin <= 194;
			36 : sin <= 198;
			37 : sin <= 202;
			38 : sin <= 206;
			39 : sin <= 209;
			40 : sin <= 213;
			41 : sin <= 216;
			42 : sin <= 220;
			43 : sin <= 223;
			44 : sin <= 226;
			45 : sin <= 229;
			46 : sin <= 231;
			47 : sin <= 234;
			48 : sin <= 237;
			49 : sin <= 239;
			50 : sin <= 241;
			51 : sin <= 243;
			52 : sin <= 245;
			53 : sin <= 247;
			54 : sin <= 248;
			55 : sin <= 250;
			56 : sin <= 251;
			57 : sin <= 252;
			58 : sin <= 253;
			59 : sin <= 254;
			60 : sin <= 255;
			61 : sin <= 255;
			62 : sin <= 256;
			63 : sin <= 256;
			64 : sin <= 256;
			65 : sin <= 256;
			66 : sin <= 256;
			67 : sin <= 255;
			68 : sin <= 255;
			69 : sin <= 254;
			70 : sin <= 253;
			71 : sin <= 252;
			72 : sin <= 251;
			73 : sin <= 250;
			74 : sin <= 248;
			75 : sin <= 247;
			76 : sin <= 245;
			77 : sin <= 243;
			78 : sin <= 241;
			79 : sin <= 239;
			80 : sin <= 237;
			81 : sin <= 234;
			82 : sin <= 231;
			83 : sin <= 229;
			84 : sin <= 226;
			85 : sin <= 223;
			86 : sin <= 220;
			87 : sin <= 216;
			88 : sin <= 213;
			89 : sin <= 209;
			90 : sin <= 206;
			91 : sin <= 202;
			92 : sin <= 198;
			93 : sin <= 194;
			94 : sin <= 190;
			95 : sin <= 185;
			96 : sin <= 181;
			97 : sin <= 177;
			98 : sin <= 172;
			99 : sin <= 167;
			100 : sin <= 162;
			101 : sin <= 157;
			102 : sin <= 152;
			103 : sin <= 147;
			104 : sin <= 142;
			105 : sin <= 137;
			106 : sin <= 132;
			107 : sin <= 126;
			108 : sin <= 121;
			109 : sin <= 115;
			110 : sin <= 109;
			111 : sin <= 104;
			112 : sin <= 98;
			113 : sin <= 92;
			114 : sin <= 86;
			115 : sin <= 80;
			116 : sin <= 74;
			117 : sin <= 68;
			118 : sin <= 62;
			119 : sin <= 56;
			120 : sin <= 50;
			121 : sin <= 44;
			122 : sin <= 38;
			123 : sin <= 31;
			124 : sin <= 25;
			125 : sin <= 19;
			126 : sin <= 13;
			127 : sin <= 6;
			128 : sin <= 0;
			129 : sin <= -6;
			130 : sin <= -13;
			131 : sin <= -19;
			132 : sin <= -25;
			133 : sin <= -31;
			134 : sin <= -38;
			135 : sin <= -44;
			136 : sin <= -50;
			137 : sin <= -56;
			138 : sin <= -62;
			139 : sin <= -68;
			140 : sin <= -74;
			141 : sin <= -80;
			142 : sin <= -86;
			143 : sin <= -92;
			144 : sin <= -98;
			145 : sin <= -104;
			146 : sin <= -109;
			147 : sin <= -115;
			148 : sin <= -121;
			149 : sin <= -126;
			150 : sin <= -132;
			151 : sin <= -137;
			152 : sin <= -142;
			153 : sin <= -147;
			154 : sin <= -152;
			155 : sin <= -157;
			156 : sin <= -162;
			157 : sin <= -167;
			158 : sin <= -172;
			159 : sin <= -177;
			160 : sin <= -181;
			161 : sin <= -185;
			162 : sin <= -190;
			163 : sin <= -194;
			164 : sin <= -198;
			165 : sin <= -202;
			166 : sin <= -206;
			167 : sin <= -209;
			168 : sin <= -213;
			169 : sin <= -216;
			170 : sin <= -220;
			171 : sin <= -223;
			172 : sin <= -226;
			173 : sin <= -229;
			174 : sin <= -231;
			175 : sin <= -234;
			176 : sin <= -237;
			177 : sin <= -239;
			178 : sin <= -241;
			179 : sin <= -243;
			180 : sin <= -245;
			181 : sin <= -247;
			182 : sin <= -248;
			183 : sin <= -250;
			184 : sin <= -251;
			185 : sin <= -252;
			186 : sin <= -253;
			187 : sin <= -254;
			188 : sin <= -255;
			189 : sin <= -255;
			190 : sin <= -256;
			191 : sin <= -256;
			192 : sin <= -256;
			193 : sin <= -256;
			194 : sin <= -256;
			195 : sin <= -255;
			196 : sin <= -255;
			197 : sin <= -254;
			198 : sin <= -253;
			199 : sin <= -252;
			200 : sin <= -251;
			201 : sin <= -250;
			202 : sin <= -248;
			203 : sin <= -247;
			204 : sin <= -245;
			205 : sin <= -243;
			206 : sin <= -241;
			207 : sin <= -239;
			208 : sin <= -237;
			209 : sin <= -234;
			210 : sin <= -231;
			211 : sin <= -229;
			212 : sin <= -226;
			213 : sin <= -223;
			214 : sin <= -220;
			215 : sin <= -216;
			216 : sin <= -213;
			217 : sin <= -209;
			218 : sin <= -206;
			219 : sin <= -202;
			220 : sin <= -198;
			221 : sin <= -194;
			222 : sin <= -190;
			223 : sin <= -185;
			224 : sin <= -181;
			225 : sin <= -177;
			226 : sin <= -172;
			227 : sin <= -167;
			228 : sin <= -162;
			229 : sin <= -157;
			230 : sin <= -152;
			231 : sin <= -147;
			232 : sin <= -142;
			233 : sin <= -137;
			234 : sin <= -132;
			235 : sin <= -126;
			236 : sin <= -121;
			237 : sin <= -115;
			238 : sin <= -109;
			239 : sin <= -104;
			240 : sin <= -98;
			241 : sin <= -92;
			242 : sin <= -86;
			243 : sin <= -80;
			244 : sin <= -74;
			245 : sin <= -68;
			246 : sin <= -62;
			247 : sin <= -56;
			248 : sin <= -50;
			249 : sin <= -44;
			250 : sin <= -38;
			251 : sin <= -31;
			252 : sin <= -25;
			253 : sin <= -19;
			254 : sin <= -13;
			255 : sin <= -6;
		endcase
		
		if(x <= 255)begin
			x <= x + 1;
		end
		else begin
			x <= 1;
			sin <= 0;
		end
	end
endmodule
	