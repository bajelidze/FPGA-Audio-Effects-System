//module delay(
//	input [31:0] sample,
//	input Enable,
//	output [15:0] left_
//);