//module tremolo_controller(
//	input 
//	);